--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   08:06:28 07/30/2017
-- Design Name:   
-- Module Name:   C:/Users/Natalia/Documents/GitHub/Assembleur/VHDL/Gates/Gates/testBench2.vhd
-- Project Name:  Gates
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: DriverGate
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY testBench2 IS
END testBench2;
 
ARCHITECTURE behavior OF testBench2 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT DriverGate
    PORT(
         x : IN  std_logic;
         F : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal x : std_logic := '0';

 	--Outputs
   signal F : std_logic;
   -- No clocks detected in port list. Replace x below with 
   -- appropriate port name 
 
   constant x_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: DriverGate PORT MAP (
          x => x,
          F => F
        );

   -- Clock process definitions
   x_process :process
   begin
		x <= '0';
		wait for x_period/2;
		x <= '1';
		wait for x_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for x_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
